module counter(input clk,output reg [3:0]q=0);

  always@(posedge clk )
    begin
        q<=q + 1;
    end
endmodule
