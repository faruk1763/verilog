module tff(input clk,rst,t,output reg q,qbar);
  always@(posedge clk or posedge rst)
    begin
    
    if(rst)
      q<=1'b0;
      else if (t)
      q<=~q;
    else
      q<=q;
      end
       assign qbar=q;
      endmodule
