module cla(
  input  g0, p0, c0,
  input  g1, p1,
  output c1, c2
);

assign c1 = g0 | (p0 & c0);
assign c2 = g1 | (p1 & g0) | (p1 & p0 & c0);

endmodule
